module ALU(
  input  [31:0] io_in1, // @[src/main/scala/npc/ALU.scala 7:16]
  input  [31:0] io_in2, // @[src/main/scala/npc/ALU.scala 7:16]
  input  [3:0]  io_op, // @[src/main/scala/npc/ALU.scala 7:16]
  output [31:0] io_out // @[src/main/scala/npc/ALU.scala 7:16]
);
  wire [31:0] add_result = io_in1 + io_in2; // @[src/main/scala/npc/ALU.scala 14:30]
  wire [31:0] sub_result = io_in1 - io_in2; // @[src/main/scala/npc/ALU.scala 15:30]
  wire [62:0] _GEN_0 = {{31'd0}, io_in1}; // @[src/main/scala/npc/ALU.scala 16:30]
  wire [62:0] sll_result = _GEN_0 << io_in2[4:0]; // @[src/main/scala/npc/ALU.scala 16:30]
  wire  slt_result = $signed(io_in1) < $signed(io_in2); // @[src/main/scala/npc/ALU.scala 17:38]
  wire  sltu_result = io_in1 < io_in2; // @[src/main/scala/npc/ALU.scala 18:32]
  wire [31:0] xor_result = io_in1 ^ io_in2; // @[src/main/scala/npc/ALU.scala 19:30]
  wire [31:0] srl_result = io_in1 >> io_in2[4:0]; // @[src/main/scala/npc/ALU.scala 20:30]
  wire [31:0] sra_result = $signed(io_in1) >>> io_in2[4:0]; // @[src/main/scala/npc/ALU.scala 21:54]
  wire [31:0] or_result = io_in1 | io_in2; // @[src/main/scala/npc/ALU.scala 22:29]
  wire [31:0] and_result = io_in1 & io_in2; // @[src/main/scala/npc/ALU.scala 23:30]
  wire [31:0] _io_out_T_1 = 4'h0 == io_op ? add_result : 32'h0; // @[src/main/scala/npc/ALU.scala 25:36]
  wire [31:0] _io_out_T_3 = 4'h1 == io_op ? sub_result : _io_out_T_1; // @[src/main/scala/npc/ALU.scala 25:36]
  wire [62:0] _io_out_T_5 = 4'h2 == io_op ? sll_result : {{31'd0}, _io_out_T_3}; // @[src/main/scala/npc/ALU.scala 25:36]
  wire [62:0] _io_out_T_7 = 4'h3 == io_op ? {{62'd0}, slt_result} : _io_out_T_5; // @[src/main/scala/npc/ALU.scala 25:36]
  wire [62:0] _io_out_T_9 = 4'h4 == io_op ? {{62'd0}, sltu_result} : _io_out_T_7; // @[src/main/scala/npc/ALU.scala 25:36]
  wire [62:0] _io_out_T_11 = 4'h5 == io_op ? {{31'd0}, xor_result} : _io_out_T_9; // @[src/main/scala/npc/ALU.scala 25:36]
  wire [62:0] _io_out_T_13 = 4'h6 == io_op ? {{31'd0}, srl_result} : _io_out_T_11; // @[src/main/scala/npc/ALU.scala 25:36]
  wire [62:0] _io_out_T_15 = 4'h7 == io_op ? {{31'd0}, sra_result} : _io_out_T_13; // @[src/main/scala/npc/ALU.scala 25:36]
  wire [62:0] _io_out_T_17 = 4'h8 == io_op ? {{31'd0}, or_result} : _io_out_T_15; // @[src/main/scala/npc/ALU.scala 25:36]
  wire [62:0] _io_out_T_19 = 4'h9 == io_op ? {{31'd0}, and_result} : _io_out_T_17; // @[src/main/scala/npc/ALU.scala 25:36]
  wire [62:0] _io_out_T_21 = 4'ha == io_op ? {{31'd0}, io_in2} : _io_out_T_19; // @[src/main/scala/npc/ALU.scala 25:36]
  assign io_out = _io_out_T_21[31:0]; // @[src/main/scala/npc/ALU.scala 25:12]
endmodule
