module LSU(
  input  [31:0] io_in_bits_aluOut, // @[src/main/scala/npc/LSU.scala 13:16]
  input  [31:0] io_in_bits_pc, // @[src/main/scala/npc/LSU.scala 13:16]
  input  [2:0]  io_in_bits_inst_type, // @[src/main/scala/npc/LSU.scala 13:16]
  input  [5:0]  io_in_bits_inst_name, // @[src/main/scala/npc/LSU.scala 13:16]
  input  [4:0]  io_in_bits_rd_addr, // @[src/main/scala/npc/LSU.scala 13:16]
  input  [10:0] io_in_bits_csr_addr, // @[src/main/scala/npc/LSU.scala 13:16]
  input  [31:0] io_in_bits_csrRdata, // @[src/main/scala/npc/LSU.scala 13:16]
  input         io_in_bits_memValid, // @[src/main/scala/npc/LSU.scala 13:16]
  input         io_in_bits_memWrite, // @[src/main/scala/npc/LSU.scala 13:16]
  input  [31:0] io_in_bits_memAddr, // @[src/main/scala/npc/LSU.scala 13:16]
  input  [31:0] io_in_bits_memWdata, // @[src/main/scala/npc/LSU.scala 13:16]
  input  [3:0]  io_in_bits_memWmask, // @[src/main/scala/npc/LSU.scala 13:16]
  input  [31:0] io_in_bits_ecall_epc, // @[src/main/scala/npc/LSU.scala 13:16]
  input  [31:0] io_in_bits_mret_epc, // @[src/main/scala/npc/LSU.scala 13:16]
  input         io_in_bits_redirect, // @[src/main/scala/npc/LSU.scala 13:16]
  input  [31:0] io_in_bits_rs1_data, // @[src/main/scala/npc/LSU.scala 13:16]
  output [31:0] io_out_bits_aluOut, // @[src/main/scala/npc/LSU.scala 13:16]
  output [31:0] io_out_bits_pc, // @[src/main/scala/npc/LSU.scala 13:16]
  output [2:0]  io_out_bits_inst_type, // @[src/main/scala/npc/LSU.scala 13:16]
  output [5:0]  io_out_bits_inst_name, // @[src/main/scala/npc/LSU.scala 13:16]
  output [4:0]  io_out_bits_rd_addr, // @[src/main/scala/npc/LSU.scala 13:16]
  output [10:0] io_out_bits_csr_addr, // @[src/main/scala/npc/LSU.scala 13:16]
  output [31:0] io_out_bits_ecall_epc, // @[src/main/scala/npc/LSU.scala 13:16]
  output [31:0] io_out_bits_mret_epc, // @[src/main/scala/npc/LSU.scala 13:16]
  output [31:0] io_out_bits_memRdata, // @[src/main/scala/npc/LSU.scala 13:16]
  output [31:0] io_out_bits_csrRdata, // @[src/main/scala/npc/LSU.scala 13:16]
  output        io_out_bits_redirect, // @[src/main/scala/npc/LSU.scala 13:16]
  output [31:0] io_out_bits_rs1_data, // @[src/main/scala/npc/LSU.scala 13:16]
  output        io_dmem_req_valid, // @[src/main/scala/npc/LSU.scala 13:16]
  output        io_dmem_req_wen, // @[src/main/scala/npc/LSU.scala 13:16]
  output [31:0] io_dmem_req_raddr, // @[src/main/scala/npc/LSU.scala 13:16]
  output [31:0] io_dmem_req_waddr, // @[src/main/scala/npc/LSU.scala 13:16]
  output [31:0] io_dmem_req_wdata, // @[src/main/scala/npc/LSU.scala 13:16]
  output [3:0]  io_dmem_req_wmask, // @[src/main/scala/npc/LSU.scala 13:16]
  input  [31:0] io_dmem_rdata // @[src/main/scala/npc/LSU.scala 13:16]
);
  assign io_out_bits_aluOut = io_in_bits_aluOut; // @[src/main/scala/npc/LSU.scala 15:17 24:23 32:28]
  assign io_out_bits_pc = io_in_bits_pc; // @[src/main/scala/npc/LSU.scala 15:17 24:23 33:24]
  assign io_out_bits_inst_type = io_in_bits_inst_type; // @[src/main/scala/npc/LSU.scala 15:17 24:23 34:31]
  assign io_out_bits_inst_name = io_in_bits_inst_name; // @[src/main/scala/npc/LSU.scala 15:17 24:23 35:31]
  assign io_out_bits_rd_addr = io_in_bits_rd_addr; // @[src/main/scala/npc/LSU.scala 15:17 24:23 39:29]
  assign io_out_bits_csr_addr = io_in_bits_csr_addr; // @[src/main/scala/npc/LSU.scala 15:17 24:23 40:30]
  assign io_out_bits_ecall_epc = io_in_bits_ecall_epc; // @[src/main/scala/npc/LSU.scala 15:17 24:23 41:31]
  assign io_out_bits_mret_epc = io_in_bits_mret_epc; // @[src/main/scala/npc/LSU.scala 15:17 24:23 42:30]
  assign io_out_bits_memRdata = io_dmem_rdata; // @[src/main/scala/npc/LSU.scala 15:17 24:23 43:30]
  assign io_out_bits_csrRdata = io_in_bits_csrRdata; // @[src/main/scala/npc/LSU.scala 15:17 24:23 44:30]
  assign io_out_bits_redirect = io_in_bits_redirect; // @[src/main/scala/npc/LSU.scala 15:17 24:23 46:30]
  assign io_out_bits_rs1_data = io_in_bits_rs1_data; // @[src/main/scala/npc/LSU.scala 15:17 24:23 38:30]
  assign io_dmem_req_valid = io_in_bits_memValid; // @[src/main/scala/npc/LSU.scala 17:23 24:23 26:27]
  assign io_dmem_req_wen = io_in_bits_memWrite; // @[src/main/scala/npc/LSU.scala 18:21 24:23 27:25]
  assign io_dmem_req_raddr = io_in_bits_memAddr; // @[src/main/scala/npc/LSU.scala 19:23 24:23 28:27]
  assign io_dmem_req_waddr = io_in_bits_memAddr; // @[src/main/scala/npc/LSU.scala 19:23 24:23 28:27]
  assign io_dmem_req_wdata = io_in_bits_memWdata; // @[src/main/scala/npc/LSU.scala 20:23 24:23 29:27]
  assign io_dmem_req_wmask = io_in_bits_memWmask; // @[src/main/scala/npc/LSU.scala 21:23 24:23 30:27]
endmodule
