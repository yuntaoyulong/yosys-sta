module EXU(
  input  [31:0] io_in_bits_imm_i, // @[src/main/scala/npc/EXU.scala 22:16]
  input  [31:0] io_in_bits_imm_s, // @[src/main/scala/npc/EXU.scala 22:16]
  input  [31:0] io_in_bits_imm_b, // @[src/main/scala/npc/EXU.scala 22:16]
  input  [31:0] io_in_bits_imm_u, // @[src/main/scala/npc/EXU.scala 22:16]
  input  [31:0] io_in_bits_imm_j, // @[src/main/scala/npc/EXU.scala 22:16]
  input  [2:0]  io_in_bits_inst_type, // @[src/main/scala/npc/EXU.scala 22:16]
  input  [5:0]  io_in_bits_inst_name, // @[src/main/scala/npc/EXU.scala 22:16]
  input  [31:0] io_in_bits_pc, // @[src/main/scala/npc/EXU.scala 22:16]
  input  [4:0]  io_in_bits_rd_addr, // @[src/main/scala/npc/EXU.scala 22:16]
  input  [10:0] io_in_bits_csr_addr, // @[src/main/scala/npc/EXU.scala 22:16]
  input  [31:0] io_in_bits_rs1_data, // @[src/main/scala/npc/EXU.scala 22:16]
  input  [31:0] io_in_bits_rs2_data, // @[src/main/scala/npc/EXU.scala 22:16]
  input  [31:0] io_in_bits_ecall_epc, // @[src/main/scala/npc/EXU.scala 22:16]
  input  [31:0] io_in_bits_mret_epc, // @[src/main/scala/npc/EXU.scala 22:16]
  input  [31:0] io_in_bits_ecall_mtvec, // @[src/main/scala/npc/EXU.scala 22:16]
  input  [31:0] io_in_bits_csr_rdata, // @[src/main/scala/npc/EXU.scala 22:16]
  output [31:0] io_out_bits_aluOut, // @[src/main/scala/npc/EXU.scala 22:16]
  output [31:0] io_out_bits_pc, // @[src/main/scala/npc/EXU.scala 22:16]
  output [2:0]  io_out_bits_inst_type, // @[src/main/scala/npc/EXU.scala 22:16]
  output [5:0]  io_out_bits_inst_name, // @[src/main/scala/npc/EXU.scala 22:16]
  output [4:0]  io_out_bits_rd_addr, // @[src/main/scala/npc/EXU.scala 22:16]
  output [10:0] io_out_bits_csr_addr, // @[src/main/scala/npc/EXU.scala 22:16]
  output [31:0] io_out_bits_csrRdata, // @[src/main/scala/npc/EXU.scala 22:16]
  output        io_out_bits_memValid, // @[src/main/scala/npc/EXU.scala 22:16]
  output        io_out_bits_memWrite, // @[src/main/scala/npc/EXU.scala 22:16]
  output [31:0] io_out_bits_memAddr, // @[src/main/scala/npc/EXU.scala 22:16]
  output [31:0] io_out_bits_memWdata, // @[src/main/scala/npc/EXU.scala 22:16]
  output [3:0]  io_out_bits_memWmask, // @[src/main/scala/npc/EXU.scala 22:16]
  output [31:0] io_out_bits_ecall_epc, // @[src/main/scala/npc/EXU.scala 22:16]
  output [31:0] io_out_bits_mret_epc, // @[src/main/scala/npc/EXU.scala 22:16]
  output        io_out_bits_redirect, // @[src/main/scala/npc/EXU.scala 22:16]
  output [31:0] io_out_bits_rs1_data // @[src/main/scala/npc/EXU.scala 22:16]
);
  wire [31:0] alu_io_in1; // @[src/main/scala/npc/EXU.scala 28:21]
  wire [31:0] alu_io_in2; // @[src/main/scala/npc/EXU.scala 28:21]
  wire [3:0] alu_io_op; // @[src/main/scala/npc/EXU.scala 28:21]
  wire [31:0] alu_io_out; // @[src/main/scala/npc/EXU.scala 28:21]
  wire  is_auipc = io_in_bits_inst_name == 6'h2d; // @[src/main/scala/npc/EXU.scala 29:41]
  wire  is_jal = io_in_bits_inst_name == 6'h2a; // @[src/main/scala/npc/EXU.scala 30:39]
  wire  is_jalr = io_in_bits_inst_name == 6'h2b; // @[src/main/scala/npc/EXU.scala 31:40]
  wire  is_beq = io_in_bits_inst_name == 6'h24; // @[src/main/scala/npc/EXU.scala 32:39]
  wire  is_bne = io_in_bits_inst_name == 6'h25; // @[src/main/scala/npc/EXU.scala 33:39]
  wire  is_blt = io_in_bits_inst_name == 6'h26; // @[src/main/scala/npc/EXU.scala 34:39]
  wire  is_bge = io_in_bits_inst_name == 6'h27; // @[src/main/scala/npc/EXU.scala 35:39]
  wire  is_bltu = io_in_bits_inst_name == 6'h28; // @[src/main/scala/npc/EXU.scala 36:40]
  wire  is_bgeu = io_in_bits_inst_name == 6'h29; // @[src/main/scala/npc/EXU.scala 37:40]
  wire  is_ecall = io_in_bits_inst_name == 6'h2f; // @[src/main/scala/npc/EXU.scala 39:41]
  wire  is_mret = io_in_bits_inst_name == 6'h32; // @[src/main/scala/npc/EXU.scala 40:40]
  wire  is_br = is_beq | is_bne | is_blt | is_bge | is_bltu | is_bgeu; // @[src/main/scala/npc/EXU.scala 47:79]
  wire [31:0] _alu_in1_T = is_auipc ? io_in_bits_pc : 32'h0; // @[src/main/scala/npc/EXU.scala 49:22]
  wire [31:0] _alu_in1_T_1 = is_br ? io_in_bits_pc : 32'h0; // @[src/main/scala/npc/EXU.scala 51:22]
  wire [31:0] _alu_in1_T_3 = is_ecall | is_mret ? io_in_bits_pc : 32'h0; // @[src/main/scala/npc/EXU.scala 52:22]
  wire  _alu_in1_T_4 = 3'h5 == io_in_bits_inst_type; // @[src/main/scala/npc/EXU.scala 48:71]
  wire [31:0] _alu_in1_T_5 = 3'h5 == io_in_bits_inst_type ? _alu_in1_T : io_in_bits_rs1_data; // @[src/main/scala/npc/EXU.scala 48:71]
  wire  _alu_in1_T_6 = 3'h6 == io_in_bits_inst_type; // @[src/main/scala/npc/EXU.scala 48:71]
  wire [31:0] _alu_in1_T_7 = 3'h6 == io_in_bits_inst_type ? io_in_bits_pc : _alu_in1_T_5; // @[src/main/scala/npc/EXU.scala 48:71]
  wire  _alu_in1_T_8 = 3'h4 == io_in_bits_inst_type; // @[src/main/scala/npc/EXU.scala 48:71]
  wire [31:0] _alu_in1_T_9 = 3'h4 == io_in_bits_inst_type ? _alu_in1_T_1 : _alu_in1_T_7; // @[src/main/scala/npc/EXU.scala 48:71]
  wire  _alu_in1_T_10 = 3'h0 == io_in_bits_inst_type; // @[src/main/scala/npc/EXU.scala 48:71]
  wire [31:0] _alu_io_in2_T = is_mret ? io_in_bits_mret_epc : 32'h0; // @[src/main/scala/npc/EXU.scala 74:14]
  wire [31:0] _alu_io_in2_T_1 = is_ecall ? io_in_bits_ecall_mtvec : _alu_io_in2_T; // @[src/main/scala/npc/EXU.scala 72:22]
  wire [31:0] _alu_io_in2_T_3 = 3'h1 == io_in_bits_inst_type ? io_in_bits_rs2_data : 32'h0; // @[src/main/scala/npc/EXU.scala 64:11]
  wire [31:0] _alu_io_in2_T_5 = 3'h2 == io_in_bits_inst_type ? io_in_bits_imm_i : _alu_io_in2_T_3; // @[src/main/scala/npc/EXU.scala 64:11]
  wire [31:0] _alu_io_in2_T_7 = 3'h3 == io_in_bits_inst_type ? io_in_bits_imm_s : _alu_io_in2_T_5; // @[src/main/scala/npc/EXU.scala 64:11]
  wire [31:0] _alu_io_in2_T_9 = _alu_in1_T_4 ? io_in_bits_imm_u : _alu_io_in2_T_7; // @[src/main/scala/npc/EXU.scala 64:11]
  wire [31:0] _alu_io_in2_T_11 = _alu_in1_T_6 ? io_in_bits_imm_j : _alu_io_in2_T_9; // @[src/main/scala/npc/EXU.scala 64:11]
  wire [31:0] _alu_io_in2_T_13 = _alu_in1_T_8 ? io_in_bits_imm_b : _alu_io_in2_T_11; // @[src/main/scala/npc/EXU.scala 64:11]
  wire [3:0] _alu_io_op_T_1 = 6'h2 == io_in_bits_inst_name ? 4'h1 : 4'h0; // @[src/main/scala/npc/EXU.scala 83:11]
  wire [3:0] _alu_io_op_T_3 = 6'h14 == io_in_bits_inst_name ? 4'h2 : _alu_io_op_T_1; // @[src/main/scala/npc/EXU.scala 83:11]
  wire [3:0] _alu_io_op_T_5 = 6'h3 == io_in_bits_inst_name ? 4'h2 : _alu_io_op_T_3; // @[src/main/scala/npc/EXU.scala 83:11]
  wire [3:0] _alu_io_op_T_7 = 6'h18 == io_in_bits_inst_name ? 4'h6 : _alu_io_op_T_5; // @[src/main/scala/npc/EXU.scala 83:11]
  wire [3:0] _alu_io_op_T_9 = 6'h7 == io_in_bits_inst_name ? 4'h6 : _alu_io_op_T_7; // @[src/main/scala/npc/EXU.scala 83:11]
  wire [3:0] _alu_io_op_T_11 = 6'h19 == io_in_bits_inst_name ? 4'h7 : _alu_io_op_T_9; // @[src/main/scala/npc/EXU.scala 83:11]
  wire [3:0] _alu_io_op_T_13 = 6'h8 == io_in_bits_inst_name ? 4'h7 : _alu_io_op_T_11; // @[src/main/scala/npc/EXU.scala 83:11]
  wire [3:0] _alu_io_op_T_15 = 6'h9 == io_in_bits_inst_name ? 4'h8 : _alu_io_op_T_13; // @[src/main/scala/npc/EXU.scala 83:11]
  wire [3:0] _alu_io_op_T_17 = 6'h1a == io_in_bits_inst_name ? 4'h8 : _alu_io_op_T_15; // @[src/main/scala/npc/EXU.scala 83:11]
  wire [3:0] _alu_io_op_T_19 = 6'h6 == io_in_bits_inst_name ? 4'h5 : _alu_io_op_T_17; // @[src/main/scala/npc/EXU.scala 83:11]
  wire [3:0] _alu_io_op_T_21 = 6'h17 == io_in_bits_inst_name ? 4'h5 : _alu_io_op_T_19; // @[src/main/scala/npc/EXU.scala 83:11]
  wire [3:0] _alu_io_op_T_23 = 6'h4 == io_in_bits_inst_name ? 4'h3 : _alu_io_op_T_21; // @[src/main/scala/npc/EXU.scala 83:11]
  wire [3:0] _alu_io_op_T_25 = 6'h15 == io_in_bits_inst_name ? 4'h3 : _alu_io_op_T_23; // @[src/main/scala/npc/EXU.scala 83:11]
  wire [3:0] _alu_io_op_T_27 = 6'h5 == io_in_bits_inst_name ? 4'h4 : _alu_io_op_T_25; // @[src/main/scala/npc/EXU.scala 83:11]
  wire [3:0] _alu_io_op_T_29 = 6'h16 == io_in_bits_inst_name ? 4'h4 : _alu_io_op_T_27; // @[src/main/scala/npc/EXU.scala 83:11]
  wire [3:0] _alu_io_op_T_31 = 6'ha == io_in_bits_inst_name ? 4'h9 : _alu_io_op_T_29; // @[src/main/scala/npc/EXU.scala 83:11]
  wire [3:0] _alu_io_op_T_33 = 6'h1b == io_in_bits_inst_name ? 4'h9 : _alu_io_op_T_31; // @[src/main/scala/npc/EXU.scala 83:11]
  wire [3:0] _alu_io_op_T_35 = 6'h2f == io_in_bits_inst_name ? 4'ha : _alu_io_op_T_33; // @[src/main/scala/npc/EXU.scala 83:11]
  wire  memRead = io_in_bits_inst_name == 6'h1c | io_in_bits_inst_name == 6'h1f | io_in_bits_inst_name == 6'h1d |
    io_in_bits_inst_name == 6'h20 | io_in_bits_inst_name == 6'h1e; // @[src/main/scala/npc/EXU.scala 114:66]
  wire  memWrite = io_in_bits_inst_name == 6'h21 | io_in_bits_inst_name == 6'h22 | io_in_bits_inst_name == 6'h23; // @[src/main/scala/npc/EXU.scala 115:68]
  wire [1:0] byteOff = alu_io_out[1:0]; // @[src/main/scala/npc/EXU.scala 116:29]
  wire [3:0] _wmask_T = 4'h1 << byteOff; // @[src/main/scala/npc/EXU.scala 123:25]
  wire [1:0] _wmask_T_1 = byteOff & 2'h2; // @[src/main/scala/npc/EXU.scala 124:37]
  wire [4:0] _wmask_T_2 = 5'h3 << _wmask_T_1; // @[src/main/scala/npc/EXU.scala 124:25]
  wire  _wmask_T_3 = 6'h21 == io_in_bits_inst_name; // @[src/main/scala/npc/EXU.scala 121:16]
  wire [3:0] _wmask_T_4 = 6'h21 == io_in_bits_inst_name ? _wmask_T : 4'h0; // @[src/main/scala/npc/EXU.scala 121:16]
  wire  _wmask_T_5 = 6'h22 == io_in_bits_inst_name; // @[src/main/scala/npc/EXU.scala 121:16]
  wire [4:0] _wmask_T_6 = 6'h22 == io_in_bits_inst_name ? _wmask_T_2 : {{1'd0}, _wmask_T_4}; // @[src/main/scala/npc/EXU.scala 121:16]
  wire [4:0] wmask = 6'h23 == io_in_bits_inst_name ? 5'hf : _wmask_T_6; // @[src/main/scala/npc/EXU.scala 121:16]
  wire [4:0] _memWdata_T_1 = {byteOff, 3'h0}; // @[src/main/scala/npc/EXU.scala 135:56]
  wire [38:0] _GEN_0 = {{31'd0}, io_in_bits_rs2_data[7:0]}; // @[src/main/scala/npc/EXU.scala 135:44]
  wire [38:0] _memWdata_T_2 = _GEN_0 << _memWdata_T_1; // @[src/main/scala/npc/EXU.scala 135:44]
  wire [4:0] _memWdata_T_5 = {_wmask_T_1, 3'h0}; // @[src/main/scala/npc/EXU.scala 136:65]
  wire [46:0] _GEN_1 = {{31'd0}, io_in_bits_rs2_data[15:0]}; // @[src/main/scala/npc/EXU.scala 136:45]
  wire [46:0] _memWdata_T_6 = _GEN_1 << _memWdata_T_5; // @[src/main/scala/npc/EXU.scala 136:45]
  wire [38:0] _memWdata_T_8 = _wmask_T_3 ? _memWdata_T_2 : {{7'd0}, io_in_bits_rs2_data}; // @[src/main/scala/npc/EXU.scala 133:27]
  wire [46:0] memWdata = _wmask_T_5 ? _memWdata_T_6 : {{8'd0}, _memWdata_T_8}; // @[src/main/scala/npc/EXU.scala 133:27]
  wire [8:0] memWmask = {4'h0,wmask}; // @[src/main/scala/npc/EXU.scala 139:23]
  wire  rs_eq = io_in_bits_rs1_data == io_in_bits_rs2_data; // @[src/main/scala/npc/EXU.scala 143:37]
  wire  rs_lt_s = $signed(io_in_bits_rs1_data) < $signed(io_in_bits_rs2_data); // @[src/main/scala/npc/EXU.scala 144:46]
  wire  rs_lt_u = io_in_bits_rs1_data < io_in_bits_rs2_data; // @[src/main/scala/npc/EXU.scala 145:39]
  wire  _do_redirect_T_1 = is_beq & rs_eq; // @[src/main/scala/npc/EXU.scala 148:17]
  wire  _do_redirect_T_2 = is_jal | is_jalr | _do_redirect_T_1; // @[src/main/scala/npc/EXU.scala 147:41]
  wire  _do_redirect_T_6 = is_blt & rs_lt_s; // @[src/main/scala/npc/EXU.scala 149:17]
  wire  _do_redirect_T_7 = _do_redirect_T_2 | is_bne & ~rs_eq | _do_redirect_T_6; // @[src/main/scala/npc/EXU.scala 148:49]
  wire  _do_redirect_T_11 = is_bltu & rs_lt_u; // @[src/main/scala/npc/EXU.scala 150:18]
  wire  _do_redirect_T_12 = _do_redirect_T_7 | is_bge & ~rs_lt_s | _do_redirect_T_11; // @[src/main/scala/npc/EXU.scala 149:53]
  wire  _do_redirect_T_16 = _do_redirect_T_12 | is_bgeu & ~rs_lt_u | is_ecall; // @[src/main/scala/npc/EXU.scala 150:55]
  ALU alu ( // @[src/main/scala/npc/EXU.scala 28:21]
    .io_in1(alu_io_in1),
    .io_in2(alu_io_in2),
    .io_op(alu_io_op),
    .io_out(alu_io_out)
  );
  assign io_out_bits_aluOut = alu_io_out; // @[src/main/scala/npc/EXU.scala 152:23 154:28 25:17]
  assign io_out_bits_pc = io_in_bits_pc; // @[src/main/scala/npc/EXU.scala 152:23 153:24 25:17]
  assign io_out_bits_inst_type = io_in_bits_inst_type; // @[src/main/scala/npc/EXU.scala 152:23 155:31 25:17]
  assign io_out_bits_inst_name = io_in_bits_inst_name; // @[src/main/scala/npc/EXU.scala 152:23 156:31 25:17]
  assign io_out_bits_rd_addr = io_in_bits_rd_addr; // @[src/main/scala/npc/EXU.scala 152:23 159:29 25:17]
  assign io_out_bits_csr_addr = io_in_bits_csr_addr; // @[src/main/scala/npc/EXU.scala 152:23 160:30 25:17]
  assign io_out_bits_csrRdata = io_in_bits_csr_rdata; // @[src/main/scala/npc/EXU.scala 152:23 167:30 25:17]
  assign io_out_bits_memValid = memRead | memWrite; // @[src/main/scala/npc/EXU.scala 129:28]
  assign io_out_bits_memWrite = io_in_bits_inst_name == 6'h21 | io_in_bits_inst_name == 6'h22 | io_in_bits_inst_name == 6'h23
    ; // @[src/main/scala/npc/EXU.scala 115:68]
  assign io_out_bits_memAddr = alu_io_out; // @[src/main/scala/npc/EXU.scala 152:23 164:29 25:17]
  assign io_out_bits_memWdata = memWdata[31:0];
  assign io_out_bits_memWmask = memWmask[3:0];
  assign io_out_bits_ecall_epc = io_in_bits_ecall_epc; // @[src/main/scala/npc/EXU.scala 152:23 168:31 25:17]
  assign io_out_bits_mret_epc = io_in_bits_mret_epc; // @[src/main/scala/npc/EXU.scala 152:23 169:30 25:17]
  assign io_out_bits_redirect = _do_redirect_T_16 | is_mret; // @[src/main/scala/npc/EXU.scala 151:18]
  assign io_out_bits_rs1_data = io_in_bits_rs1_data; // @[src/main/scala/npc/EXU.scala 152:23 161:30 25:17]
  assign alu_io_in1 = 3'h0 == io_in_bits_inst_type ? _alu_in1_T_3 : _alu_in1_T_9; // @[src/main/scala/npc/EXU.scala 48:71]
  assign alu_io_in2 = _alu_in1_T_10 ? _alu_io_in2_T_1 : _alu_io_in2_T_13; // @[src/main/scala/npc/EXU.scala 64:11]
  assign alu_io_op = 6'h32 == io_in_bits_inst_name ? 4'ha : _alu_io_op_T_35; // @[src/main/scala/npc/EXU.scala 83:11]
endmodule
