// module EbreakDetector(
//   input io_ebreak
// );
//   import "DPI-C" function void ebreak_handler();
  
//   always @(posedge io_ebreak) begin
//     ebreak_handler();
//   end

  
// endmodule