module WBU(
  input  [31:0] io_in_bits_aluOut, // @[src/main/scala/npc/WBU.scala 17:16]
  input  [31:0] io_in_bits_pc, // @[src/main/scala/npc/WBU.scala 17:16]
  input  [2:0]  io_in_bits_inst_type, // @[src/main/scala/npc/WBU.scala 17:16]
  input  [5:0]  io_in_bits_inst_name, // @[src/main/scala/npc/WBU.scala 17:16]
  input  [4:0]  io_in_bits_rd_addr, // @[src/main/scala/npc/WBU.scala 17:16]
  input  [10:0] io_in_bits_csr_addr, // @[src/main/scala/npc/WBU.scala 17:16]
  input  [31:0] io_in_bits_ecall_epc, // @[src/main/scala/npc/WBU.scala 17:16]
  input  [31:0] io_in_bits_mret_epc, // @[src/main/scala/npc/WBU.scala 17:16]
  input  [31:0] io_in_bits_memRdata, // @[src/main/scala/npc/WBU.scala 17:16]
  input  [31:0] io_in_bits_csrRdata, // @[src/main/scala/npc/WBU.scala 17:16]
  input         io_in_bits_redirect, // @[src/main/scala/npc/WBU.scala 17:16]
  input  [31:0] io_in_bits_rs1_data, // @[src/main/scala/npc/WBU.scala 17:16]
  output [4:0]  io_rfout_rd_addr, // @[src/main/scala/npc/WBU.scala 17:16]
  output [31:0] io_rfout_rd_data, // @[src/main/scala/npc/WBU.scala 17:16]
  output        io_rfout_rd_wen, // @[src/main/scala/npc/WBU.scala 17:16]
  output [10:0] io_rfout_csr_addr, // @[src/main/scala/npc/WBU.scala 17:16]
  output [31:0] io_rfout_csr_wdata, // @[src/main/scala/npc/WBU.scala 17:16]
  output        io_rfout_csr_wen, // @[src/main/scala/npc/WBU.scala 17:16]
  output        io_rfout_do_ecall, // @[src/main/scala/npc/WBU.scala 17:16]
  output [31:0] io_rfout_ecall_epc, // @[src/main/scala/npc/WBU.scala 17:16]
  output        io_rfout_do_mret, // @[src/main/scala/npc/WBU.scala 17:16]
  input         io_out_ready, // @[src/main/scala/npc/WBU.scala 17:16]
  output [31:0] io_out_bits_dnpc, // @[src/main/scala/npc/WBU.scala 17:16]
  output        io_out_bits_redirect // @[src/main/scala/npc/WBU.scala 17:16]
);
  wire [31:0] pc4 = io_in_bits_pc + 32'h4; // @[src/main/scala/npc/WBU.scala 19:29]
  wire [1:0] byteOff = io_in_bits_aluOut[1:0]; // @[src/main/scala/npc/WBU.scala 22:36]
  wire [4:0] _b_T = {byteOff, 3'h0}; // @[src/main/scala/npc/WBU.scala 23:46]
  wire [31:0] _b_T_1 = io_in_bits_memRdata >> _b_T; // @[src/main/scala/npc/WBU.scala 23:34]
  wire [7:0] b = _b_T_1[7:0]; // @[src/main/scala/npc/WBU.scala 23:52]
  wire [4:0] _h_T_1 = {io_in_bits_aluOut[1], 4'h0}; // @[src/main/scala/npc/WBU.scala 24:59]
  wire [31:0] _h_T_2 = io_in_bits_memRdata >> _h_T_1; // @[src/main/scala/npc/WBU.scala 24:34]
  wire [15:0] h = _h_T_2[15:0]; // @[src/main/scala/npc/WBU.scala 24:65]
  wire [23:0] _loadData_T_1 = b[7] ? 24'hffffff : 24'h0; // @[src/main/scala/npc/WBU.scala 27:28]
  wire [31:0] _loadData_T_2 = {_loadData_T_1,b}; // @[src/main/scala/npc/WBU.scala 27:23]
  wire [31:0] _loadData_T_4 = {24'h0,b}; // @[src/main/scala/npc/WBU.scala 28:24]
  wire [15:0] _loadData_T_6 = h[15] ? 16'hffff : 16'h0; // @[src/main/scala/npc/WBU.scala 29:28]
  wire [31:0] _loadData_T_7 = {_loadData_T_6,h}; // @[src/main/scala/npc/WBU.scala 29:23]
  wire [31:0] _loadData_T_9 = {16'h0,h}; // @[src/main/scala/npc/WBU.scala 30:24]
  wire  _loadData_T_10 = 6'h1c == io_in_bits_inst_name; // @[src/main/scala/npc/WBU.scala 25:72]
  wire [31:0] _loadData_T_11 = 6'h1c == io_in_bits_inst_name ? _loadData_T_2 : io_in_bits_memRdata; // @[src/main/scala/npc/WBU.scala 25:72]
  wire  _loadData_T_12 = 6'h1f == io_in_bits_inst_name; // @[src/main/scala/npc/WBU.scala 25:72]
  wire [31:0] _loadData_T_13 = 6'h1f == io_in_bits_inst_name ? _loadData_T_4 : _loadData_T_11; // @[src/main/scala/npc/WBU.scala 25:72]
  wire  _loadData_T_14 = 6'h1d == io_in_bits_inst_name; // @[src/main/scala/npc/WBU.scala 25:72]
  wire [31:0] _loadData_T_15 = 6'h1d == io_in_bits_inst_name ? _loadData_T_7 : _loadData_T_13; // @[src/main/scala/npc/WBU.scala 25:72]
  wire  _loadData_T_16 = 6'h20 == io_in_bits_inst_name; // @[src/main/scala/npc/WBU.scala 25:72]
  wire [31:0] _loadData_T_17 = 6'h20 == io_in_bits_inst_name ? _loadData_T_9 : _loadData_T_15; // @[src/main/scala/npc/WBU.scala 25:72]
  wire  _loadData_T_18 = 6'h1e == io_in_bits_inst_name; // @[src/main/scala/npc/WBU.scala 25:72]
  wire [31:0] loadData = 6'h1e == io_in_bits_inst_name ? io_in_bits_memRdata : _loadData_T_17; // @[src/main/scala/npc/WBU.scala 25:72]
  wire [31:0] _wbData_T_1 = _loadData_T_10 ? loadData : io_in_bits_aluOut; // @[src/main/scala/npc/WBU.scala 36:68]
  wire [31:0] _wbData_T_3 = _loadData_T_12 ? loadData : _wbData_T_1; // @[src/main/scala/npc/WBU.scala 36:68]
  wire [31:0] _wbData_T_5 = _loadData_T_14 ? loadData : _wbData_T_3; // @[src/main/scala/npc/WBU.scala 36:68]
  wire [31:0] _wbData_T_7 = _loadData_T_16 ? loadData : _wbData_T_5; // @[src/main/scala/npc/WBU.scala 36:68]
  wire [31:0] _wbData_T_9 = _loadData_T_18 ? loadData : _wbData_T_7; // @[src/main/scala/npc/WBU.scala 36:68]
  wire [31:0] _wbData_T_11 = 6'h2a == io_in_bits_inst_name ? pc4 : _wbData_T_9; // @[src/main/scala/npc/WBU.scala 36:68]
  wire [31:0] _wbData_T_13 = 6'h2b == io_in_bits_inst_name ? pc4 : _wbData_T_11; // @[src/main/scala/npc/WBU.scala 36:68]
  wire [31:0] _wbData_T_15 = 6'h31 == io_in_bits_inst_name ? io_in_bits_csrRdata : _wbData_T_13; // @[src/main/scala/npc/WBU.scala 36:68]
  wire [31:0] _wbData_T_17 = 6'h30 == io_in_bits_inst_name ? io_in_bits_csrRdata : _wbData_T_15; // @[src/main/scala/npc/WBU.scala 36:68]
  wire [31:0] _wbData_T_19 = 6'h2f == io_in_bits_inst_name ? io_in_bits_ecall_epc : _wbData_T_17; // @[src/main/scala/npc/WBU.scala 36:68]
  wire  _io_rfout_rd_wen_T_3 = io_in_bits_inst_type != 3'h0; // @[src/main/scala/npc/WBU.scala 64:35]
  wire  _io_rfout_csr_wen_T_1 = io_in_bits_inst_name == 6'h30; // @[src/main/scala/npc/WBU.scala 67:92]
  wire [31:0] _io_rfout_csr_wdata_T_1 = io_in_bits_csrRdata | io_in_bits_rs1_data; // @[src/main/scala/npc/WBU.scala 71:31]
  assign io_rfout_rd_addr = io_in_bits_rd_addr; // @[src/main/scala/npc/WBU.scala 53:14 57:23 58:26]
  assign io_rfout_rd_data = 6'h32 == io_in_bits_inst_name ? io_in_bits_mret_epc : _wbData_T_19; // @[src/main/scala/npc/WBU.scala 36:68]
  assign io_rfout_rd_wen = io_in_bits_inst_type != 3'h3 & io_in_bits_inst_type != 3'h4 & _io_rfout_rd_wen_T_3; // @[src/main/scala/npc/WBU.scala 63:99]
  assign io_rfout_csr_addr = io_in_bits_csr_addr; // @[src/main/scala/npc/WBU.scala 53:14 57:23 59:27]
  assign io_rfout_csr_wdata = _io_rfout_csr_wen_T_1 ? io_in_bits_rs1_data : _io_rfout_csr_wdata_T_1; // @[src/main/scala/npc/WBU.scala 68:34]
  assign io_rfout_csr_wen = io_in_bits_inst_name == 6'h31 | io_in_bits_inst_name == 6'h30; // @[src/main/scala/npc/WBU.scala 67:67]
  assign io_rfout_do_ecall = io_in_bits_inst_name == 6'h2f; // @[src/main/scala/npc/WBU.scala 74:45]
  assign io_rfout_ecall_epc = io_in_bits_pc; // @[src/main/scala/npc/WBU.scala 53:14 57:23 80:28]
  assign io_rfout_do_mret = io_in_bits_inst_name == 6'h32; // @[src/main/scala/npc/WBU.scala 75:44]
  assign io_out_bits_dnpc = io_in_bits_aluOut; // @[src/main/scala/npc/WBU.scala 54:22]
  assign io_out_bits_redirect = io_in_bits_redirect; // @[src/main/scala/npc/WBU.scala 55:26]
endmodule
